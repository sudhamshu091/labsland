module mux_2_to_1();
